GENERATOR
$time=0 a=0 b=1 sum=0 carry=0
DRIVER
$time=0 a=0 b=1 sum=0 carry=0
MONITOR
$time=1 a=0 b=1 sum=1 carry=0
SCOREBOARD
$time=1 a=0 b=1 sum=1 carry=0
Correct
___________________
GENERATOR
$time=1 a=1 b=1 sum=0 carry=0
DRIVER
$time=1 a=1 b=1 sum=0 carry=0
MONITOR
$time=7 a=1 b=1 sum=0 carry=1
SCOREBOARD
$time=7 a=1 b=1 sum=0 carry=1
Correct
___________________
GENERATOR
$time=7 a=0 b=1 sum=0 carry=0
DRIVER
$time=7 a=0 b=1 sum=0 carry=0
MONITOR
$time=13 a=0 b=1 sum=1 carry=0
SCOREBOARD
$time=13 a=0 b=1 sum=1 carry=0
Correct
___________________
GENERATOR
$time=13 a=0 b=1 sum=0 carry=0
DRIVER
$time=13 a=0 b=1 sum=0 carry=0
MONITOR
$time=19 a=0 b=1 sum=1 carry=0
SCOREBOARD
$time=19 a=0 b=1 sum=1 carry=0
Correct
___________________
GENERATOR
$time=19 a=1 b=1 sum=0 carry=0
DRIVER
$time=19 a=1 b=1 sum=0 carry=0
MONITOR
$time=25 a=1 b=1 sum=0 carry=1
SCOREBOARD
$time=25 a=1 b=1 sum=0 carry=1
Correct
___________________
GENERATOR
$time=25 a=1 b=1 sum=0 carry=0
DRIVER
$time=25 a=1 b=1 sum=0 carry=0
MONITOR
$time=31 a=1 b=1 sum=0 carry=1
SCOREBOARD
$time=31 a=1 b=1 sum=0 carry=1
Correct
___________________
GENERATOR
$time=31 a=1 b=1 sum=0 carry=0
DRIVER
$time=31 a=1 b=1 sum=0 carry=0
MONITOR
$time=37 a=1 b=1 sum=0 carry=1
SCOREBOARD
$time=37 a=1 b=1 sum=0 carry=1
Correct
___________________
GENERATOR
$time=37 a=1 b=1 sum=0 carry=0
DRIVER
$time=37 a=1 b=1 sum=0 carry=0
MONITOR
$time=43 a=1 b=1 sum=0 carry=1
SCOREBOARD
$time=43 a=1 b=1 sum=0 carry=1
Correct
___________________
GENERATOR
$time=43 a=0 b=1 sum=0 carry=0
DRIVER
$time=43 a=0 b=1 sum=0 carry=0
MONITOR
$time=49 a=0 b=1 sum=1 carry=0
SCOREBOARD
$time=49 a=0 b=1 sum=1 carry=0
Correct
___________________
GENERATOR
$time=49 a=1 b=1 sum=0 carry=0
DRIVER
$time=49 a=1 b=1 sum=0 carry=0
MONITOR
$time=55 a=1 b=1 sum=0 carry=1
SCOREBOARD
$time=55 a=1 b=1 sum=0 carry=1
Correct
___________________
GENERATOR
$time=55 a=0 b=1 sum=0 carry=0
DRIVER
$time=55 a=0 b=1 sum=0 carry=0
MONITOR
$time=61 a=0 b=1 sum=1 carry=0
SCOREBOARD
$time=61 a=0 b=1 sum=1 carry=0
Correct
___________________
GENERATOR
$time=61 a=0 b=0 sum=0 carry=0
DRIVER
$time=61 a=0 b=0 sum=0 carry=0
MONITOR
$time=67 a=0 b=0 sum=0 carry=0
SCOREBOARD
$time=67 a=0 b=0 sum=0 carry=0
Correct
___________________
GENERATOR
$time=67 a=1 b=1 sum=0 carry=0
DRIVER
$time=67 a=1 b=1 sum=0 carry=0
MONITOR
$time=73 a=1 b=1 sum=0 carry=1
SCOREBOARD
$time=73 a=1 b=1 sum=0 carry=1
Correct
___________________
GENERATOR
$time=73 a=0 b=0 sum=0 carry=0
DRIVER
$time=73 a=0 b=0 sum=0 carry=0
MONITOR
$time=79 a=0 b=0 sum=0 carry=0
SCOREBOARD
$time=79 a=0 b=0 sum=0 carry=0
Correct
___________________
GENERATOR
$time=79 a=0 b=1 sum=0 carry=0
DRIVER
$time=79 a=0 b=1 sum=0 carry=0
MONITOR
$time=85 a=0 b=1 sum=1 carry=0
SCOREBOARD
$time=85 a=0 b=1 sum=1 carry=0
Correct
___________________
GENERATOR
$time=85 a=1 b=1 sum=0 carry=0
DRIVER
$time=85 a=1 b=1 sum=0 carry=0
MONITOR
$time=91 a=1 b=1 sum=0 carry=1
SCOREBOARD
$time=91 a=1 b=1 sum=0 carry=1
Correct
___________________
GENERATOR
$time=91 a=0 b=0 sum=0 carry=0
DRIVER
$time=91 a=0 b=0 sum=0 carry=0
MONITOR
$time=97 a=0 b=0 sum=0 carry=0
SCOREBOARD
$time=97 a=0 b=0 sum=0 carry=0
Correct
___________________
GENERATOR
$time=97 a=1 b=1 sum=0 carry=0
DRIVER
$time=97 a=1 b=1 sum=0 carry=0
MONITOR
$time=103 a=1 b=1 sum=0 carry=1
SCOREBOARD
$time=103 a=1 b=1 sum=0 carry=1
Correct
___________________
GENERATOR
$time=103 a=0 b=0 sum=0 carry=0
DRIVER
$time=103 a=0 b=0 sum=0 carry=0
MONITOR
$time=109 a=0 b=0 sum=0 carry=0
SCOREBOARD
$time=109 a=0 b=0 sum=0 carry=0
Correct
___________________
GENERATOR
$time=109 a=1 b=0 sum=0 carry=0
DRIVER
$time=109 a=1 b=0 sum=0 carry=0
MONITOR
$time=115 a=1 b=0 sum=1 carry=0
SCOREBOARD
$time=115 a=1 b=0 sum=1 carry=0
Correct
___________________
$finish at simulation time                  120
           V C S   S i m u l a t i o n   R e p o r t 
