interface interf;
  
    logic d0;
    logic d1;
    logic s;
    logic y;
    endinterface
    
