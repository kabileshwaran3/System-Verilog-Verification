interface inter;
  logic clk;
  logic rst;
  logic [7:0]data_in;
  logic enable;
  logic [2:0]addrs;
  logic [7:0]data_out;
  
endinterface
         
