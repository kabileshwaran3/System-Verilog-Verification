interface interf;
  logic [3:0]a,b;
  logic cin;
  logic [3:0]sum;
  logic cout;
endinterface
