Memory Created
Time Delay                   0
start randomize value 
                   0  a=0,b=1, cin=1, sum=0, carry=0
value Assigned
driver class
                   0  a=0,b=1, cin=1, sum=0, carry=0
Value passed to interface
monitor block
                   2  a=0,b=1, cin=1, sum=0, carry=1
Full adder opertion
scoreboard signal
                   2  a=0,b=1, cin=1, sum=0, carry=1
Expected output = Original output
correct
Memory Created
Time Delay                   3
start randomize value 
                   3  a=1,b=0, cin=0, sum=0, carry=0
value Assigned
driver class
                   3  a=1,b=0, cin=0, sum=0, carry=0
Value passed to interface
monitor block
                   5  a=1,b=0, cin=0, sum=1, carry=0
Full adder opertion
scoreboard signal
                   5  a=1,b=0, cin=0, sum=1, carry=0
Expected output = Original output
correct
Memory Created
Time Delay                   6
start randomize value 
                   6  a=0,b=0, cin=1, sum=0, carry=0
value Assigned
driver class
                   6  a=0,b=0, cin=1, sum=0, carry=0
Value passed to interface
monitor block
                   8  a=0,b=0, cin=1, sum=1, carry=0
Full adder opertion
scoreboard signal
                   8  a=0,b=0, cin=1, sum=1, carry=0
Expected output = Original output
correct
Memory Created
Time Delay                   9
start randomize value 
                   9  a=1,b=0, cin=0, sum=0, carry=0
value Assigned
driver class
                   9  a=1,b=0, cin=0, sum=0, carry=0
Value passed to interface
monitor block
                  11  a=1,b=0, cin=0, sum=1, carry=0
Full adder opertion
scoreboard signal
                  11  a=1,b=0, cin=0, sum=1, carry=0
Expected output = Original output
correct
Memory Created
Time Delay                  12
start randomize value 
                  12  a=0,b=1, cin=0, sum=0, carry=0
value Assigned
driver class
                  12  a=0,b=1, cin=0, sum=0, carry=0
Value passed to interface
monitor block
                  14  a=0,b=1, cin=0, sum=1, carry=0
Full adder opertion
scoreboard signal
                  14  a=0,b=1, cin=0, sum=1, carry=0
Expected output = Original output
correct
$finish at simulation time                   15
           V C S   S i m u l a t i o n   R e p o r t 
