xcelium> run
Generator Class
*****start randomize value *********
                   0  a=1101,b=1111, cin=1, sum=0000, cout=0
driver class
*****######## Enter into driver class #########*********
                   0  a=1101,b=1111, cin=1, sum=0000, cout=0
Value passed to interface
########## Enter into monitor block ########
*****monitor block*********
                   3  a=1101,b=1111, cin=1, sum=1101, cout=1
Ripple Carry adder opertion
*****scoreboard signal*********
                   3  a=1101,b=1111, cin=1, sum=1101, cout=1
Scoreboard: Correct output
Generator Class
*****start randomize value *********
                   3  a=0001,b=1110, cin=0, sum=0000, cout=0
driver class
*****######## Enter into driver class #########*********
                   3  a=0001,b=1110, cin=0, sum=0000, cout=0
Value passed to interface
########## Enter into monitor block ########
*****monitor block*********
                   7  a=0001,b=1110, cin=0, sum=1111, cout=0
Ripple Carry adder opertion
*****scoreboard signal*********
                   7  a=0001,b=1110, cin=0, sum=1111, cout=0
Scoreboard: Correct output
Generator Class
*****start randomize value *********
                   7  a=1100,b=1001, cin=0, sum=0000, cout=0
driver class
*****######## Enter into driver class #########*********
                   7  a=1100,b=1001, cin=0, sum=0000, cout=0
Value passed to interface
########## Enter into monitor block ########
*****monitor block*********
                  11  a=1100,b=1001, cin=0, sum=0101, cout=1
Ripple Carry adder opertion
*****scoreboard signal*********
                  11  a=1100,b=1001, cin=0, sum=0101, cout=1
Scoreboard: Correct output
Generator Class
*****start randomize value *********
                  11  a=1110,b=1001, cin=0, sum=0000, cout=0
driver class
*****######## Enter into driver class #########*********
                  11  a=1110,b=1001, cin=0, sum=0000, cout=0
Value passed to interface
########## Enter into monitor block ########
*****monitor block*********
                  15  a=1110,b=1001, cin=0, sum=0111, cout=1
Ripple Carry adder opertion
*****scoreboard signal*********
                  15  a=1110,b=1001, cin=0, sum=0111, cout=1
Scoreboard: Correct output
Generator Class
*****start randomize value *********
                  15  a=0101,b=0101, cin=0, sum=0000, cout=0
driver class
*****######## Enter into driver class #########*********
                  15  a=0101,b=0101, cin=0, sum=0000, cout=0
Value passed to interface
########## Enter into monitor block ########
*****monitor block*********
                  19  a=0101,b=0101, cin=0, sum=1010, cout=0
Ripple Carry adder opertion
*****scoreboard signal*********
                  19  a=0101,b=0101, cin=0, sum=1010, cout=0
Scoreboard: Correct output
Generator Class
*****start randomize value *********
                  19  a=0010,b=1100, cin=0, sum=0000, cout=0
driver class
*****######## Enter into driver class #########*********
                  19  a=0010,b=1100, cin=0, sum=0000, cout=0
Value passed to interface
########## Enter into monitor block ########
*****monitor block*********
                  23  a=0010,b=1100, cin=0, sum=1110, cout=0
Ripple Carry adder opertion
*****scoreboard signal*********
                  23  a=0010,b=1100, cin=0, sum=1110, cout=0
Scoreboard: Correct output
Generator Class
*****start randomize value *********
                  23  a=1001,b=1110, cin=1, sum=0000, cout=0
driver class
*****######## Enter into driver class #########*********
                  23  a=1001,b=1110, cin=1, sum=0000, cout=0
Value passed to interface
########## Enter into monitor block ########
*****monitor block*********
                  27  a=1001,b=1110, cin=1, sum=1000, cout=1
Ripple Carry adder opertion
*****scoreboard signal*********
                  27  a=1001,b=1110, cin=1, sum=1000, cout=1
Scoreboard: Correct output
Generator Class
*****start randomize value *********
                  27  a=1010,b=1000, cin=0, sum=0000, cout=0
driver class
*****######## Enter into driver class #########*********
                  27  a=1010,b=1000, cin=0, sum=0000, cout=0
Value passed to interface
########## Enter into monitor block ########
*****monitor block*********
                  31  a=1010,b=1000, cin=0, sum=0010, cout=1
Ripple Carry adder opertion
*****scoreboard signal*********
                  31  a=1010,b=1000, cin=0, sum=0010, cout=1
Scoreboard: Correct output
Generator Class
*****start randomize value *********
                  31  a=0000,b=0101, cin=0, sum=0000, cout=0
driver class
*****######## Enter into driver class #########*********
                  31  a=0000,b=0101, cin=0, sum=0000, cout=0
Value passed to interface
########## Enter into monitor block ########
*****monitor block*********
                  35  a=0000,b=0101, cin=0, sum=0101, cout=0
Ripple Carry adder opertion
*****scoreboard signal*********
                  35  a=0000,b=0101, cin=0, sum=0101, cout=0
Scoreboard: Correct output
Generator Class
*****start randomize value *********
                  35  a=0110,b=0010, cin=0, sum=0000, cout=0
driver class
*****######## Enter into driver class #########*********
                  35  a=0110,b=0010, cin=0, sum=0000, cout=0
Value passed to interface
########## Enter into monitor block ########
*****monitor block*********
                  39  a=0110,b=0010, cin=0, sum=1000, cout=0
Ripple Carry adder opertion
*****scoreboard signal*********
                  39  a=0110,b=0010, cin=0, sum=1000, cout=0
Scoreboard: Correct output
