interface inter();
  logic clk,rst;
  logic mode;
  logic [3:0]count;
endinterface
